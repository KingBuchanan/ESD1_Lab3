--
-- YOUR HEADER GOES HERE
--
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.std_logic_unsigned.ALL;
ENTITY raminfr IS
  PORT (
    clk : IN std_logic;
    reset_n : IN std_logic;
    we_n : IN std_logic;
    be_n : IN std_logic_vector(3 DOWNTO 0);
    addr : IN std_logic_vector(11 DOWNTO 0);
    din : IN std_logic_vector(31 DOWNTO 0);
    dout : OUT std_logic_vector(31 DOWNTO 0)
);
END ENTITY raminfr;

ARCHITECTURE rtl OF raminfr IS
  TYPE ram_type_1 IS ARRAY (4095 DOWNTO 0) OF std_logic_vector (7 DOWNTO 0);
  TYPE ram_type_2 IS ARRAY (4095 DOWNTO 0) OF std_logic_vector (7 DOWNTO 0);
  TYPE ram_type_3 IS ARRAY (4095 DOWNTO 0) OF std_logic_vector (7 DOWNTO 0);
  TYPE ram_type_4 IS ARRAY (4095 DOWNTO 0) OF std_logic_vector (7 DOWNTO 0);
  SIGNAL RAM : ram_type_1;
  SIGNAL RAM_2 : ram_type_2;
  SIGNAL RAM_3 : ram_type_3;
  SIGNAL RAM_4 : ram_type_4;
  SIGNAL read_addr : std_logic_vector(11 DOWNTO 0);
BEGIN
  RamBlock : PROCESS(clk) BEGIN
    IF (clk'event AND clk = '1') THEN
      IF (reset_n = '0') THEN
        read_addr <= (OTHERS => '0');
      ELSIF (we_n = '0')&(be_n='0000') THEN
        RAM(conv_integer(addr)) <= din(31 downto 23);
        RAM_2(conv_integer(addr)) <= din(23 downto 15);
        RAM_3(conv_integer(addr)) <= din(15 downto 7);
        RAM_4(conv_integer(addr)) <= din(7 downto 0);
      END IF;
      read_addr <= addr;
    END IF;
  END PROCESS RamBlock;
  dout <= (RAM & RAM_2 & RAM_3 &RAM_4)(conv_integer(read_addr));
END ARCHITECTURE rtl;